module caculate_exp_thapphan(thapphan,so_mu)