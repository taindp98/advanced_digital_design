`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: VHT
// Engineer: taindp@viettel.com.vn
// 
// Create Date: 24/05/2019 02:56:40 PM
// Design Name: 
// Module Name: find_1_first.v
// Project Name: KTSNC 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module find_1_first(I,position,flag);
      input       [24:0]I;
      output	flag;
      output	[4:0]position;

      wire [4:0]  position1;
      
      assign	flag=~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]
                      &~I[16]&~I[15]&~I[14]&~I[13]&~I[12]&~I[11]&~I[10]&~I[9]
      		    &~I[8]&~I[7]&~I[6]&~I[5]&~I[4]&~I[3]&~I[2]&~I[1]&~I[0];

      assign 	position1[0]=(~I[24]&I[23])
                              |(~I[24]&~I[22]&I[21])
                              |(~I[24]&~I[22]&~I[20]&I[19])
      	                  |(~I[24]&~I[22]&~I[20]&~I[18]&I[17])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&I[15])
                               |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&I[13])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&I[11])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&I[9])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&I[7])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&~I[6]&I[5])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&~I[6]&~I[4]&I[3])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&~I[6]&~I[4]&~I[2]&I[1]);

      assign	position1[1]=(~I[24]&~I[23]&I[22])
                              |(~I[24]&~I[23]&I[21])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&I[18])
                              |(~I[24]&~I[23]&~I[20]&~I[19]&I[17])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&I[14])
                              |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&I[13])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&I[10])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&I[9])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&I[6])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&I[5])
                              |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&~I[4]&~I[3]&I[2])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&~I[4]&~I[3]&I[1]);

      assign	position1[2]=(~I[24]&~I[23]&~I[22]&~I[21]&I[20])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&I[19])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&I[18])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&I[17])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[12])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[11])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[10])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[9])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[4])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[3])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[2]) 
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[1]);

      assign	position1[3]=(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[16])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[15])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[14])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[13])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[12])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[11])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[10])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[9])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&~I[8]&~I[7]&~I[6]&~I[5]&~I[4]&~I[3]&~I[2]&~I[1]&I[0]);

      assign	position1[4]=(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&~I[16]&~I[15]
                        &~I[14]&~I[13]&~I[12]&~I[11]&~I[10]&~I[9])&(I[8]|I[7]|I[6]|I[5]|I[4]|I[3]|I[2]|I[1]|I[0]);
      assign      position=flag?5'b00000:position1;

endmodule
