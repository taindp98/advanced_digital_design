module AU_FLOATING_POINT_TESTBENCH;
	reg [31:0] A,B;
	reg [1:0]sel;

	wire [31:0]result;
	wire underflag,overflag;

	AU_FLOATING_POINT uut(A,B,sel,overflag,underflag,result);

	initial begin
////////////////////////////////


		A=32'h00000000;
		B=32'h00000000;
		sel=2'b00;
	#100
		A=32'h00000000;
		B=32'h00000000;
		sel=2'b01;
	#100
		A=32'h00000000;
		B=32'h00000000;
		sel=2'b10;
	#100
		A=32'h00000000;
		B=32'h00000000;
		sel=2'b11;
	#100
//////////////////////////////////////
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b00;
		#100
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b01;
		#100
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b10;
		#100
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b11;
		#100
/////////////////////////////////////////\
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b00;
		#100
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b01;
		#100
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b10;
		#100
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b11;
		#100
//////////////////////////////////////////////
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b00;
		#100
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b01;
		#100
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b10;
		#100
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b11;
		#100	
////////////////////////////////////////////////////
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b00;
		#100
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b01;
		#100
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b10;
		#100
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b11;
		#100
		
//////////////////////////////////////////////////////////
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b00;
		#100
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b01;
		#100
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b10;
		#100
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b11;
		#100
///////////////////////////////////////////////////////////
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b11;
	end

endmodule
