`timescale 1ns / 1ns
module multiplier_tb;
   wire [31:0]result;
    wire underflag,overflag;

    reg [31:0]A,B;
  


    multiplier uut(.A(A),
                .B(B),
                .overflag(overflag),
                .underflag(underflag),
                .result(result));


    initial
        begin
            A = 32'b00111110000000000000000000000000; //0.125
            B = 32'b01000001000101100000000000000000; //9.375
    
            #50

////////////////////////////////////////////////////////////////////////////////
            A = 32'b10111110000000000000000000000000; //-0.125
            B = 32'b11000001000101100000000000000000; //-9.375
      
            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b10111110000000000000000000000000; //-0.125
            B = 32'b11000001000101100000000000000000; //-9.375
  
            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b00000000000000000000000000000000; //0
            B = 32'b11000001000101100000000000000000; //-9.375
      
            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b01111111100000000000000000000000; //+vo cung
            B = 32'b11000001000101100000000000000000; //-9.375
      
            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b01111111100000000000000000000000; //+vo cung
            B = 32'b11111111100000000000000000000000; //-vo cung
         
            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b01111111100000000000000000000000; //+vo cung
            B = 32'b01111111100000000000000000000000; //+vo cung
         

            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b00111000010100011011011100010111; //0.00005
            B = 32'b01100000101011010111100011101100; //10^20
    

            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b00111000010100011011011100010111; //0.00005
            B = 32'b01100111010100111100001000011100; //10^25

            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b00000000000000000000000000000000; //0
            B = 32'b01111111100000000000000000000000; //+vo cung
      
        
            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b00000000000000000000000000000000; //0
            B = 32'b11111111100000000000000000000000; //-vo cung

            #50
//////////////////////////////////////////////////////////////////////////////////
            A = 32'b00111000010100011011011100010111; //0.00005
            B = 32'b01100111010100111100001000011100; //10^25
      

        end
endmodule
