`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: VHT
// Engineer: taindp@viettel.com.vn
// 
// Create Date: 24/05/2019 02:56:40 PM
// Design Name: 
// Module Name: add_sub_tb.v
// Project Name: KTSNC 
// Target Devices: 
// Tool Versions: 
// Description: testbench add_sub
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module add_sub_tb;
	wire	[31:0]result;
	wire underflow,overflow;

	reg [31:0]A,B;
	reg	add_or_sub;


	add_sub uut(.A(A),
				.B(B),
				.add_or_sub(add_or_sub),
				.overflow(overflow),
				.underflow(underflow),
				.result(result));


	initial
		begin
			A = 32'b00111110000000000000000000000000; //0.125
			B = 32'b01000001000101100000000000000000; //9.375
			add_or_sub = 0;
							//rs=9.5 // 01000001000110000000000000000000
			#50
///////////////////////////////////////////////////////////////////////////////////
			A = 32'b00111110000000000000000000000000; //0.125
			B = 32'b01000001000101100000000000000000; //9.375
			add_or_sub = 1;
					//result=-9.25   //11000001000101000000000000000000
			#50
////////////////////////////////////////////////////////////////////////////////
			A = 32'b10111110000000000000000000000000; //-0.125
			B = 32'b11000001000101100000000000000000; //-9.375
			add_or_sub = 0;
					//result=-9.5  
			#50
//////////////////////////////////////////////////////////////////////////////////
			A = 32'b10111110000000000000000000000000; //-0.125
			B = 32'b11000001000101100000000000000000; //-9.375
			add_or_sub = 1;
					//result=9.25
			#50
//////////////////////////////////////////////////////////////////////////////////
			A = 32'b00000000000000000000000000000000; //0
			B = 32'b11000001000101100000000000000000; //-9.375
			add_or_sub = 1;
					//result=9.375
			#50
//////////////////////////////////////////////////////////////////////////////////
			A = 32'b01111111100000000000000000000000; //+vo cung
			B = 32'b11000001000101100000000000000000; //-9.375
			add_or_sub = 1;
					//result=Inf
			#50
//////////////////////////////////////////////////////////////////////////////////
			A = 32'b01111111100000000000000000000000; //+vo cung
			B = 32'b11111111100000000000000000000000; //-vo cung
			add_or_sub = 1;
					//result=Inf
			#50
//////////////////////////////////////////////////////////////////////////////////
			A = 32'b01111111100000000000000000000000; //+vo cung
			B = 32'b01111111100000000000000000000000; //+vo cung
			add_or_sub = 1;
					//result=NaN

			#50
//////////////////////////////////////////////////////////////////////////////////
			A = 32'b00111000010100011011011100010111; //0.00005
			B = 32'b01100000101011010111100011101100; //10^20
			add_or_sub = 0;
					//

			#50
//////////////////////////////////////////////////////////////////////////////////
			A = 32'b00111000010100011011011100010111; //0.00005
			B = 32'b01100111010100111100001000011100; //10^24
			add_or_sub = 1;
					//
			#50;
		end
endmodule
