module AU_FLOATING_POINT_TESTBENCH;
	reg [31:0] A,B;
	reg [1:0]sel;

	wire [31:0]result;
	wire underflag,overflag;

	AU_FLOATING_POINT uut(A,B,sel,overflag,underflag,result);

	initial begin
////////////////////////////////


		A=32'h00000000;
		B=32'h00000000;
		sel=2'b00;
	#100
		A=32'h00000000;
		B=32'h00000000;
		sel=2'b01;
	#100
		A=32'h00000000;
		B=32'h00000000;
		sel=2'b10;
	#100
		A=32'h00000000;
		B=32'h00000000;
		sel=2'b11;
	#100
//////////////////////////////////////
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b00;
		#100
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b01;
		#100
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b10;
		#100
		A=32'h00000000;
		B=32'hFF800000;
		sel=2'b11;
		#100
/////////////////////////////////////////\
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b00;
		#100
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b01;
		#100
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b10;
		#100
		A=32'hFF800000;
		B=32'h7F800000;
		sel=2'b11;
		#100
//////////////////////////////////////////////
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b00;
		#100
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b01;
		#100
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b10;
		#100
		A=32'hFF800000;
		B=32'h00000000;
		sel=2'b11;
		#100	
////////////////////////////////////////////////////
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b00;
		#100
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b01;
		#100
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b10;
		#100
		A=32'h44fc6000; //2019
		B=32'hc4f9e000; //-1999
		sel=2'b11;
		#100
		
//////////////////////////////////////////////////////////
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b00;
		#100
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b01;
		#100
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b10;
		#100
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b11;
		#100

		A=32'b01001100000000000000000000000000; //2^25
		B=32'b01000000000000000000000000000000 ; //2
		sel=2'b01;

		#100

		B=32'b01001100000000000000000000000000; //2^25
		A=32'b01000000000000000000000000000000 ; //2
		sel=2'b01;

		#100
		A=32'hc05f5c29;
		B=32'b01000010110010010000111101011100;
		sel=2'b10;

		#100
		A=32'hc4b772e1;
		B=32'h3f2dd2f2;
		sel=2'b10;

		#100
		A=32'h3dfbe76d;
		B=32'h3f2d9168;
		sel=2'b10;

		#100
		A=32'b01111011111000000000000000000000;
		B=32'b01110001110101000000000000000000;
		sel=2'b10;


	#100
///////////////////////////////////////////////////////////
		A=32'hc4fc6fae;
		B=32'h3f449ba6;
		sel=2'b11;
	end

endmodule
